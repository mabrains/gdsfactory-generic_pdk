** test_straight_heater_doped_strip circuit for GenericPDK
* ========================================================================
* SPDX-FileCopyrightText: 2023 Mabrains Company
* Licensed under the GNU GENERAL PUBLIC License, Version 3.0 (the "License");
* you may not use this file except in compliance with the License.
*
*                    GNU GENERAL PUBLIC LICENSE
*                       Version 3, 29 June 2007
*
* This program is free software: you can redistribute it and/or modify
* it under the terms of the GNU General Public License as published
* by the Free Software Foundation, either 3 of the License, or
* (at your option) any later version.
* 
* This program is distributed in the hope that it will be useful,
* but WITHOUT ANY WARRANTY; without even the implied warranty of
* MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
* GNU General Public License for more details.
* 
* You should have received a copy of the GNU General Public License
* along with this program.  If not, see <https://www.gnu.org/licenses/>.
* SPDX-License-Identifier: GPL-3.0
* ========================================================================

.subckt test_straight_heater_doped_strip pin1 pin2 hp_pin hn_pin
*.PININFO pin1:B pin2:B hp_pin:B hn_pin:B
Pheater1 pin1 net1 hn_pin hp_pin straight_heater_doped_strip length=320.0 nsections=3
+ heater_width=2.0 heater_gap=0.8 via_stack_gap=0.0 width=0.5 xoffset_tip1=0.2 xoffset_tip2=0.4
Pheater2 net1 net2 hn_pin hp_pin straight_heater_doped_strip length=320.0 nsections=3
+ heater_width=2.0 heater_gap=0.8 via_stack_gap=0.0 width=0.5 xoffset_tip1=0.2 xoffset_tip2=0.4
Pheater3 net2 net3 hn_pin hp_pin straight_heater_doped_strip length=320.0 nsections=3
+ heater_width=2.0 heater_gap=0.8 via_stack_gap=0.0 width=0.5 xoffset_tip1=0.2 xoffset_tip2=0.4
Pheater4 net3 net4 hn_pin hp_pin straight_heater_doped_strip length=320.0 nsections=3
+ heater_width=2.0 heater_gap=0.8 via_stack_gap=0.0 width=0.5 xoffset_tip1=0.2 xoffset_tip2=0.4
Pheater5 net4 pin2 hn_pin hp_pin straight_heater_doped_strip length=320.0 nsections=3
+ heater_width=2.0 heater_gap=0.8 via_stack_gap=0.0 width=0.5 xoffset_tip1=0.2 xoffset_tip2=0.4
.ends
.end
