** test_mmi1x2_with_sbend circuit for GenericPDK
* ========================================================================
* SPDX-FileCopyrightText: 2023 Mabrains Company
* Licensed under the GNU GENERAL PUBLIC License, Version 3.0 (the "License");
* you may not use this file except in compliance with the License.
*
*                    GNU GENERAL PUBLIC LICENSE
*                       Version 3, 29 June 2007
*
* This program is free software: you can redistribute it and/or modify
* it under the terms of the GNU General Public License as published
* by the Free Software Foundation, either 3 of the License, or
* (at your option) any later version.
* 
* This program is distributed in the hope that it will be useful,
* but WITHOUT ANY WARRANTY; without even the implied warranty of
* MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
* GNU General Public License for more details.
* 
* You should have received a copy of the GNU General Public License
* along with this program.  If not, see <https://www.gnu.org/licenses/>.
* SPDX-License-Identifier: GPL-3.0
* ========================================================================

.subckt test_mmi1x2_with_sbend pin1 pin3 pin2
*.PININFO pin1:B pin3:B pin2:B
Pmmi1 pin2 net5 net6 mmi1x2_with_sbend
Pmmi2 net1 net6 net5 mmi1x2_with_sbend
Pmmi3 pin1 net2 net1 mmi1x2_with_sbend
Pmmi4 net2 net3 net4 mmi1x2_with_sbend
Pmmi5 pin3 net4 net3 mmi1x2_with_sbend
.ends
.end
