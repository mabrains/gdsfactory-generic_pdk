** test_ring_single_pn circuit for GenericPDK
* ========================================================================
* SPDX-FileCopyrightText: 2023 Mabrains Company
* Licensed under the GNU GENERAL PUBLIC License, Version 3.0 (the "License");
* you may not use this file except in compliance with the License.
*
*                    GNU GENERAL PUBLIC LICENSE
*                       Version 3, 29 June 2007
*
* This program is free software: you can redistribute it and/or modify
* it under the terms of the GNU General Public License as published
* by the Free Software Foundation, either 3 of the License, or
* (at your option) any later version.
* 
* This program is distributed in the hope that it will be useful,
* but WITHOUT ANY WARRANTY; without even the implied warranty of
* MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
* GNU General Public License for more details.
* 
* You should have received a copy of the GNU General Public License
* along with this program.  If not, see <https://www.gnu.org/licenses/>.
* SPDX-License-Identifier: GPL-3.0
* ========================================================================

.subckt test_ring_single_pn pin1 pin2
*.PININFO pin1:B pin2:B
Pring1 pin1 net4 ring_single_pn gap=0.3 radius=5.0 doping_angle=250 length_x=0.1 length_y=0.1
Pring2 net4 net1 ring_single_pn gap=0.3 radius=5.0 doping_angle=250 length_x=0.1 length_y=0.1
Pring3 net1 net2 ring_single_pn gap=0.3 radius=5.0 doping_angle=250 length_x=0.1 length_y=0.1
Pring4 net3 net2 ring_single_pn gap=0.3 radius=5.0 doping_angle=250 length_x=0.1 length_y=0.1
Pring5 net3 pin2 ring_single_pn gap=0.3 radius=5.0 doping_angle=250 length_x=0.1 length_y=0.1
.ends
.end
