** test_ring_single circuit for GenericPDK
* ========================================================================
* SPDX-FileCopyrightText: 2023 Mabrains Company
* Licensed under the GNU GENERAL PUBLIC License, Version 3.0 (the "License");
* you may not use this file except in compliance with the License.
*
*                    GNU GENERAL PUBLIC LICENSE
*                       Version 3, 29 June 2007
*
* This program is free software: you can redistribute it and/or modify
* it under the terms of the GNU General Public License as published
* by the Free Software Foundation, either 3 of the License, or
* (at your option) any later version.
* 
* This program is distributed in the hope that it will be useful,
* but WITHOUT ANY WARRANTY; without even the implied warranty of
* MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
* GNU General Public License for more details.
* 
* You should have received a copy of the GNU General Public License
* along with this program.  If not, see <https://www.gnu.org/licenses/>.
* SPDX-License-Identifier: GPL-3.0
* ========================================================================

.subckt test_ring_single pin1 pin2
*.iopin pin1
*.iopin pin2
Pring1 pin1 net4 ring_single gap=0.2 radius=10.0 length_x=4.0 length_y=0.6
Pring2 net4 net1 ring_single gap=0.2 radius=10.0 length_x=4.0 length_y=0.6
Pring3 net1 net2 ring_single gap=0.2 radius=10.0 length_x=4.0 length_y=0.6
Pring4 net3 net2 ring_single gap=0.2 radius=10.0 length_x=4.0 length_y=0.6
Pring5 net3 pin2 ring_single gap=0.2 radius=10.0 length_x=4.0 length_y=0.6
.ends
.end
