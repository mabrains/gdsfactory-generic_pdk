** test_mzi2x2_2x2_phase_shifter circuit for GenericPDK
* ========================================================================
* SPDX-FileCopyrightText: 2023 Mabrains Company
* Licensed under the GNU GENERAL PUBLIC License, Version 3.0 (the "License");
* you may not use this file except in compliance with the License.
*
*                    GNU GENERAL PUBLIC LICENSE
*                       Version 3, 29 June 2007
*
* This program is free software: you can redistribute it and/or modify
* it under the terms of the GNU General Public License as published
* by the Free Software Foundation, either 3 of the License, or
* (at your option) any later version.
* 
* This program is distributed in the hope that it will be useful,
* but WITHOUT ANY WARRANTY; without even the implied warranty of
* MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
* GNU General Public License for more details.
* 
* You should have received a copy of the GNU General Public License
* along with this program.  If not, see <https://www.gnu.org/licenses/>.
* SPDX-License-Identifier: GPL-3.0
* ========================================================================

.subckt test_mzi2x2_2x2_phase_shifter pin2 pin3 pin1 pin4
*.PININFO pin2:B pin3:B pin1:B pin4:B
Pmzi1 pin1 net3 net4 pin2 mzi2x2_2x2_phase_shifter delta_length=10.0 length_y=2.0 length_x=0.1
Pmzi2 net3 net5 net6 net4 mzi2x2_2x2_phase_shifter delta_length=10.0 length_y=2.0 length_x=0.1
Pmzi3 net6 net1 net2 net6 mzi2x2_2x2_phase_shifter delta_length=10.0 length_y=2.0 length_x=0.1
Pmzi4 net1 pin3 pin4 net2 mzi2x2_2x2_phase_shifter delta_length=10.0 length_y=2.0 length_x=0.1
.ends
.end
