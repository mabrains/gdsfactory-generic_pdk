** test_mzm circuit for GenericPDK
* ========================================================================
* SPDX-FileCopyrightText: 2023 Mabrains Company
* Licensed under the GNU GENERAL PUBLIC License, Version 3.0 (the "License");
* you may not use this file except in compliance with the License.
*
*                    GNU GENERAL PUBLIC LICENSE
*                       Version 3, 29 June 2007
*
* This program is free software: you can redistribute it and/or modify
* it under the terms of the GNU General Public License as published
* by the Free Software Foundation, either 3 of the License, or
* (at your option) any later version.
* 
* This program is distributed in the hope that it will be useful,
* but WITHOUT ANY WARRANTY; without even the implied warranty of
* MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
* GNU General Public License for more details.
* 
* You should have received a copy of the GNU General Public License
* along with this program.  If not, see <https://www.gnu.org/licenses/>.
* SPDX-License-Identifier: GPL-3.0
* ========================================================================

.subckt test_mzm pin2 pin1 pin3
*.PININFO pin2:B pin1:B pin3:B
Pmzm1 net1 net2 mzm length_x=500 length_y=2.0 delta_length=0.0
Pmzm2 net2 net3 mzm length_x=500 length_y=2.0 delta_length=0.0
Pmzm3 pin1 net3 mzm length_x=500 length_y=2.0 delta_length=0.0
Pmzm4 net3 net4 mzm length_x=500 length_y=2.0 delta_length=0.0
Pmzm5 net4 pin3 mzm length_x=500 length_y=2.0 delta_length=0.0
.ends
.end
