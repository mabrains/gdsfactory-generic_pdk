** test_mzit circuit for GenericPDK
* ========================================================================
* SPDX-FileCopyrightText: 2023 Mabrains Company
* Licensed under the GNU GENERAL PUBLIC License, Version 3.0 (the "License");
* you may not use this file except in compliance with the License.
*
*                    GNU GENERAL PUBLIC LICENSE
*                       Version 3, 29 June 2007
*
* This program is free software: you can redistribute it and/or modify
* it under the terms of the GNU General Public License as published
* by the Free Software Foundation, either 3 of the License, or
* (at your option) any later version.
* 
* This program is distributed in the hope that it will be useful,
* but WITHOUT ANY WARRANTY; without even the implied warranty of
* MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
* GNU General Public License for more details.
* 
* You should have received a copy of the GNU General Public License
* along with this program.  If not, see <https://www.gnu.org/licenses/>.
* SPDX-License-Identifier: GPL-3.0
* ========================================================================

.subckt test_mzit pin2 pin1 pin4 pin3
*.PININFO pin2:B pin1:B pin4:B pin3:B
Pmzi1 pin1 pin2 net3 net4 mzit w0=0.5 w1=0.45 w2=0.55 dy=2.0 delta_length=10.0 length=1.0
+ coupler_length1=5.0 coupler_length2=10.0 coupler_gap1=0.2 coupler_gap2=0.3 taper_length=5.0
Pmzi2 net6 net5 net4 net3 mzit w0=0.5 w1=0.45 w2=0.55 dy=2.0 delta_length=10.0 length=1.0
+ coupler_length1=5.0 coupler_length2=10.0 coupler_gap1=0.2 coupler_gap2=0.3 taper_length=5.0
Pmzi3 net6 net5 net2 net1 mzit w0=0.5 w1=0.45 w2=0.55 dy=2.0 delta_length=10.0 length=1.0
+ coupler_length1=5.0 coupler_length2=10.0 coupler_gap1=0.2 coupler_gap2=0.3 taper_length=5.0
Pmzi4 net2 net1 pin4 pin3 mzit w0=0.5 w1=0.45 w2=0.55 dy=2.0 delta_length=10.0 length=1.0
+ coupler_length1=5.0 coupler_length2=10.0 coupler_gap1=0.2 coupler_gap2=0.3 taper_length=5.0
.ends
.end
