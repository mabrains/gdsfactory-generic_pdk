** test_mmi2x2 circuit for GenericPDK
* ========================================================================
* SPDX-FileCopyrightText: 2023 Mabrains Company
* Licensed under the GNU GENERAL PUBLIC License, Version 3.0 (the "License");
* you may not use this file except in compliance with the License.
*
*                    GNU GENERAL PUBLIC LICENSE
*                       Version 3, 29 June 2007
*
* This program is free software: you can redistribute it and/or modify
* it under the terms of the GNU General Public License as published
* by the Free Software Foundation, either 3 of the License, or
* (at your option) any later version.
* 
* This program is distributed in the hope that it will be useful,
* but WITHOUT ANY WARRANTY; without even the implied warranty of
* MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
* GNU General Public License for more details.
* 
* You should have received a copy of the GNU General Public License
* along with this program.  If not, see <https://www.gnu.org/licenses/>.
* SPDX-License-Identifier: GPL-3.0
* ========================================================================

.subckt test_mmi2x2 pin1 pin2 pin3 pin4
*.PININFO pin1:B pin2:B pin3:B pin4:B
Pmmi2 pin2 pin1 net1 net2 mmi2x2 width=0.5 width_taper=1 length_taper=10 length_mmi=5.5
+ width_mmi=2.5 gap_mmi=0.25
Pmmi1 net2 net1 net3 net4 mmi2x2 width=0.5 width_taper=1 length_taper=10 length_mmi=5.5
+ width_mmi=2.5 gap_mmi=0.25
Pmmi3 net4 net3 net6 net5 mmi2x2 width=0.5 width_taper=1 length_taper=10 length_mmi=5.5
+ width_mmi=2.5 gap_mmi=0.25
Pmmi4 net5 net6 pin3 pin4 mmi2x2 width=0.5 width_taper=1 length_taper=10 length_mmi=5.5
+ width_mmi=2.5 gap_mmi=0.25
.ends
.end
